CONSTANT  SHL  :  std_logic_vector(4 downto 0)  := "00000";
CONSTANT  SHR  :  std_logic_vector(4 downto 0)  := "00001";
CONSTANT  ADD  :  std_logic_vector(4 downto 0)  := "00010";--first bit must be 0 and sub is the opposite (also in inc and dec)
CONSTANT  SUB  :  std_logic_vector(4 downto 0)  := "00011";
CONSTANT  RLC  :  std_logic_vector(4 downto 0)  := "00100";
CONSTANT  RRC  :  std_logic_vector(4 downto 0)  := "00101";
CONSTANT  myAND  :  std_logic_vector(4 downto 0)  := "00110";
CONSTANT  myOR  :  std_logic_vector(4 downto 0)  := "00111";
CONSTANT  INC  :  std_logic_vector(4 downto 0)  := "01000";
CONSTANT  DEC  :  std_logic_vector(4 downto 0)  :=  "01001";
CONSTANT  SETC  :  std_logic_vector(4 downto 0)  := "01010";
CONSTANT  CLC  :  std_logic_vector(4 downto 0)  := "01011";
CONSTANT  myNOT  :  std_logic_vector(4 downto 0)  := "01100";
CONSTANT  NEG  :  std_logic_vector(4 downto 0)  := "01101";
CONSTANT  STD  :  std_logic_vector(4 downto 0)  := "01110";
CONSTANT  MOV  :  std_logic_vector(4 downto 0)  := "01111";
CONSTANT  LDM  :  std_logic_vector(4 downto 0)  := "10000";
CONSTANT  LDD  :  std_logic_vector(4 downto 0)  := "10001";